library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;

-- running on board: Cyclone 5 GX Starter Kit 

entity SevenSegmentDriver is	
	port (
		data:     in STD_LOGIC_VECTOR(3 downto 0);
		en:       in STD_LOGIC;
		q:       out STD_LOGIC_VECTOR (6 downto 0)
	);	
end entity;


architecture immediate of SevenSegmentDriver is
begin		
	process (data,en)		
	begin	
	   if en='0' then
		   q <= "1111111";
		else
		   case data is 
			when "0000" =>     -- 0
			    q(0) <= '0';
			    q(1) <= '0';
			    q(2) <= '0';
			    q(3) <= '0';
			    q(4) <= '0';
			    q(5) <= '0';
			    q(6) <= '1';
		   when "0001" =>   -- 1
			    q(0) <= '1';
			    q(1) <= '0';
			    q(2) <= '0';
			    q(3) <= '1';
			    q(4) <= '1';
			    q(5) <= '1';
			    q(6) <= '1';
		   when "0010" =>  -- 2
			    q(0) <= '0';
			    q(1) <= '0';
			    q(2) <= '1';
			    q(3) <= '0';
			    q(4) <= '0';
			    q(5) <= '1';
			    q(6) <= '0';
		   when "0011"  =>  -- 3
			    q(0) <= '0';
			    q(1) <= '0';
			    q(2) <= '0';
			    q(3) <= '0';
			    q(4) <= '1';
			    q(5) <= '1';
			    q(6) <= '0';
		   when "0100"  =>  -- 4
			    q(0) <= '1';
			    q(1) <= '0';
			    q(2) <= '0';
			    q(3) <= '1';
			    q(4) <= '1';
			    q(5) <= '0';
			    q(6) <= '0';
		   when "0101" => -- 5
			    q(0) <= '0';
			    q(1) <= '1';
			    q(2) <= '0';
			    q(3) <= '0';
			    q(4) <= '1';
			    q(5) <= '0';
			    q(6) <= '0';
		   when "0110" => -- 6
			    q(0) <= '0';
			    q(1) <= '1';
			    q(2) <= '0';
			    q(3) <= '0';
			    q(4) <= '0';
			    q(5) <= '0';
			    q(6) <= '0';
		   when "0111" =>  -- 7
			    q(0) <= '0';
			    q(1) <= '0';
			    q(2) <= '0';
			    q(3) <= '1';
			    q(4) <= '1';
			    q(5) <= '1';
			    q(6) <= '1';
		   when "1000" =>  -- 8
			    q(0) <= '0';
			    q(1) <= '0';
			    q(2) <= '0';
			    q(3) <= '0';
			    q(4) <= '0';
			    q(5) <= '0';
			    q(6) <= '0';
		   when "1001"  =>  -- 9
			    q(0) <= '0';
			    q(1) <= '0';
			    q(2) <= '0';
			    q(3) <= '0';
			    q(4) <= '1';
			    q(5) <= '0';
			    q(6) <= '0';
		   when "1010"  =>  -- A
			    q(0) <= '0';
			    q(1) <= '0';
			    q(2) <= '0';
			    q(3) <= '1';
			    q(4) <= '0';
			    q(5) <= '0';
			    q(6) <= '0';
		   when "1011"  =>  -- b
			    q(0) <= '1';
			    q(1) <= '1';
			    q(2) <= '0';
			    q(3) <= '0';
			    q(4) <= '0';
			    q(5) <= '0';
			    q(6) <= '0';
		   when "1100"  => -- C
			    q(0) <= '0';
			    q(1) <= '1';
			    q(2) <= '1';
			    q(3) <= '0';
			    q(4) <= '0';
			    q(5) <= '0';
			    q(6) <= '1';
		   when "1101"  =>  -- d
			    q(0) <= '1';
			    q(1) <= '0';
			    q(2) <= '0';
			    q(3) <= '0';
			    q(4) <= '0';
			    q(5) <= '1';
			    q(6) <= '0';
		   when "1110"  =>  -- E
			    q(0) <= '0';
			    q(1) <= '1';
			    q(2) <= '1';
			    q(3) <= '0';
			    q(4) <= '0';
			    q(5) <= '0';
			    q(6) <= '0';
		   when "1111" =>  -- F
			    q(0) <= '0';
			    q(1) <= '1';
			    q(2) <= '1';
			    q(3) <= '1';
			    q(4) <= '0';
			    q(5) <= '0';
			    q(6) <= '0';
         end case;
		end if;
	end process;	
	
end immediate;


